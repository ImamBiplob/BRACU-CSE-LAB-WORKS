module problem1_18301276 (y,a,b,c);
	input a,b,c;
	output y;
	
	assign y = ~(~(~(a&a)&~(b&b)&c)&~(~(a&a)&b&~(c&c))&~(a&~(b&b)&~(c&c))&~(a&b&c));
endmodule